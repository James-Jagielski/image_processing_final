magic
tech sky130A
timestamp 1695693994
<< nwell >>
rect -135 1340 205 2165
<< nmos >>
rect -65 1165 -50 1265
rect -25 1165 -10 1265
rect 40 1165 70 1265
rect 120 1165 135 1265
rect -65 675 -50 775
rect -25 675 -10 775
rect 40 675 70 775
rect 120 675 135 775
<< pmos >>
rect -65 1890 -50 1990
rect 0 1890 15 1990
rect 65 1890 80 1990
rect 120 1890 135 1990
rect -65 1360 -50 1460
rect 0 1360 15 1460
rect 65 1360 80 1460
rect 120 1360 135 1460
<< ndiff >>
rect -115 1250 -65 1265
rect -115 1180 -100 1250
rect -80 1180 -65 1250
rect -115 1165 -65 1180
rect -50 1165 -25 1265
rect -10 1250 40 1265
rect -10 1180 5 1250
rect 25 1180 40 1250
rect -10 1165 40 1180
rect 70 1250 120 1265
rect 70 1180 85 1250
rect 105 1180 120 1250
rect 70 1165 120 1180
rect 135 1250 185 1265
rect 135 1180 150 1250
rect 170 1180 185 1250
rect 135 1165 185 1180
rect -115 760 -65 775
rect -115 690 -100 760
rect -80 690 -65 760
rect -115 675 -65 690
rect -50 675 -25 775
rect -10 760 40 775
rect -10 690 5 760
rect 25 690 40 760
rect -10 675 40 690
rect 70 760 120 775
rect 70 690 85 760
rect 105 690 120 760
rect 70 675 120 690
rect 135 760 185 775
rect 135 690 150 760
rect 170 690 185 760
rect 135 675 185 690
<< pdiff >>
rect -115 1975 -65 1990
rect -115 1905 -100 1975
rect -80 1905 -65 1975
rect -115 1890 -65 1905
rect -50 1975 0 1990
rect -50 1905 -35 1975
rect -15 1905 0 1975
rect -50 1890 0 1905
rect 15 1975 65 1990
rect 15 1905 30 1975
rect 50 1905 65 1975
rect 15 1890 65 1905
rect 80 1890 120 1990
rect 135 1975 185 1990
rect 135 1905 150 1975
rect 170 1905 185 1975
rect 135 1890 185 1905
rect -115 1445 -65 1460
rect -115 1375 -100 1445
rect -80 1375 -65 1445
rect -115 1360 -65 1375
rect -50 1445 0 1460
rect -50 1375 -35 1445
rect -15 1375 0 1445
rect -50 1360 0 1375
rect 15 1445 65 1460
rect 15 1375 30 1445
rect 50 1375 65 1445
rect 15 1360 65 1375
rect 80 1360 120 1460
rect 135 1445 185 1460
rect 135 1375 150 1445
rect 170 1375 185 1445
rect 135 1360 185 1375
<< ndiffc >>
rect -100 1180 -80 1250
rect 5 1180 25 1250
rect 85 1180 105 1250
rect 150 1180 170 1250
rect -100 690 -80 760
rect 5 690 25 760
rect 85 690 105 760
rect 150 690 170 760
<< pdiffc >>
rect -100 1905 -80 1975
rect -35 1905 -15 1975
rect 30 1905 50 1975
rect 150 1905 170 1975
rect -100 1375 -80 1445
rect -35 1375 -15 1445
rect 30 1375 50 1445
rect 150 1375 170 1445
<< psubdiff >>
rect -40 630 10 645
rect -40 560 -25 630
rect -5 560 10 630
rect -40 545 10 560
rect 95 630 145 645
rect 95 560 110 630
rect 130 560 145 630
rect 95 545 145 560
<< nsubdiff >>
rect -60 2130 -10 2145
rect -60 2060 -45 2130
rect -25 2060 -10 2130
rect -60 2045 -10 2060
rect 80 2130 130 2145
rect 80 2060 95 2130
rect 115 2060 130 2130
rect 80 2045 130 2060
<< psubdiffcont >>
rect -25 560 -5 630
rect 110 560 130 630
<< nsubdiffcont >>
rect -45 2060 -25 2130
rect 95 2060 115 2130
<< poly >>
rect -65 1990 -50 2005
rect 0 1990 15 2005
rect 65 1990 80 2005
rect 120 1990 135 2005
rect -65 1460 -50 1890
rect 0 1625 15 1890
rect -25 1615 15 1625
rect -25 1595 -15 1615
rect 5 1595 15 1615
rect -25 1585 15 1595
rect -25 1550 15 1560
rect -25 1530 -15 1550
rect 5 1530 15 1550
rect -25 1520 15 1530
rect 0 1460 15 1520
rect 65 1460 80 1890
rect 120 1830 135 1890
rect 105 1820 145 1830
rect 105 1800 115 1820
rect 135 1800 145 1820
rect 105 1790 145 1800
rect 105 1755 145 1765
rect 105 1735 115 1755
rect 135 1735 145 1755
rect 105 1725 145 1735
rect 120 1460 135 1725
rect -65 1265 -50 1360
rect 0 1345 15 1360
rect 65 1345 80 1360
rect -25 1330 15 1345
rect 55 1330 80 1345
rect -25 1265 -10 1330
rect 55 1280 70 1330
rect 40 1265 70 1280
rect 120 1265 135 1360
rect -65 775 -50 1165
rect -25 1110 -10 1165
rect -25 1100 15 1110
rect -25 1080 -15 1100
rect 5 1080 15 1100
rect -25 1070 15 1080
rect -25 1035 15 1045
rect -25 1015 -15 1035
rect 5 1015 15 1035
rect -25 1005 15 1015
rect -25 775 -10 1005
rect 40 775 70 1165
rect 120 1000 135 1165
rect 120 985 155 1000
rect 140 955 155 985
rect 115 945 155 955
rect 115 925 125 945
rect 145 925 155 945
rect 115 915 155 925
rect 95 865 135 875
rect 95 845 105 865
rect 125 845 135 865
rect 95 835 135 845
rect 120 775 135 835
rect -65 530 -50 675
rect -25 660 -10 675
rect 40 530 70 675
rect 120 660 135 675
rect -90 520 -50 530
rect -90 500 -80 520
rect -60 500 -50 520
rect -90 490 -50 500
rect 30 520 70 530
rect 30 500 40 520
rect 60 500 70 520
rect 30 490 70 500
<< polycont >>
rect -15 1595 5 1615
rect -15 1530 5 1550
rect 115 1800 135 1820
rect 115 1735 135 1755
rect -15 1080 5 1100
rect -15 1015 5 1035
rect 125 925 145 945
rect 105 845 125 865
rect -80 500 -60 520
rect 40 500 60 520
<< locali >>
rect -55 2130 -15 2140
rect -55 2060 -45 2130
rect -25 2060 -15 2130
rect -55 2050 -15 2060
rect 85 2130 125 2140
rect 85 2060 95 2130
rect 115 2060 125 2130
rect 85 2050 125 2060
rect -110 1975 -70 1985
rect -110 1905 -100 1975
rect -80 1905 -70 1975
rect -110 1895 -70 1905
rect -45 1975 -5 1985
rect -45 1905 -35 1975
rect -15 1905 -5 1975
rect -45 1895 -5 1905
rect 20 1975 60 1985
rect 20 1905 30 1975
rect 50 1905 60 1975
rect 20 1895 60 1905
rect 140 1975 180 1985
rect 140 1905 150 1975
rect 170 1905 180 1975
rect 140 1895 180 1905
rect -25 1665 -5 1895
rect 140 1870 160 1895
rect 65 1850 160 1870
rect 65 1765 85 1850
rect 105 1820 145 1830
rect 105 1800 115 1820
rect 135 1810 145 1820
rect 135 1800 185 1810
rect 105 1790 185 1800
rect 65 1755 145 1765
rect 65 1745 115 1755
rect 105 1735 115 1745
rect 135 1735 145 1755
rect 105 1725 145 1735
rect 165 1705 185 1790
rect 140 1685 185 1705
rect -25 1645 55 1665
rect -25 1615 15 1625
rect -25 1605 -15 1615
rect -65 1595 -15 1605
rect 5 1595 15 1615
rect -65 1585 15 1595
rect -65 1500 -45 1585
rect 35 1560 55 1645
rect -25 1550 55 1560
rect -25 1530 -15 1550
rect 5 1540 55 1550
rect 5 1530 15 1540
rect -25 1520 15 1530
rect -65 1480 -25 1500
rect -45 1455 -25 1480
rect 140 1455 160 1685
rect -110 1445 -70 1455
rect -110 1375 -100 1445
rect -80 1375 -70 1445
rect -110 1365 -70 1375
rect -45 1445 -5 1455
rect -45 1375 -35 1445
rect -15 1375 -5 1445
rect -45 1365 -5 1375
rect 20 1445 60 1455
rect 20 1375 30 1445
rect 50 1375 60 1445
rect 20 1365 60 1375
rect 140 1445 180 1455
rect 140 1375 150 1445
rect 170 1375 180 1445
rect 140 1365 180 1375
rect -25 1305 -5 1365
rect 140 1340 160 1365
rect 95 1320 160 1340
rect -25 1285 35 1305
rect 15 1260 35 1285
rect 95 1260 115 1320
rect -110 1250 -70 1260
rect -110 1180 -100 1250
rect -80 1180 -70 1250
rect -110 1170 -70 1180
rect -5 1250 35 1260
rect -5 1180 5 1250
rect 25 1180 35 1250
rect -5 1170 35 1180
rect 15 1150 35 1170
rect 75 1250 115 1260
rect 75 1180 85 1250
rect 105 1180 115 1250
rect 75 1170 115 1180
rect 140 1250 180 1260
rect 140 1180 150 1250
rect 170 1180 180 1250
rect 140 1170 180 1180
rect 15 1130 55 1150
rect -25 1100 15 1110
rect -25 1090 -15 1100
rect -65 1080 -15 1090
rect 5 1080 15 1100
rect -65 1070 15 1080
rect -65 985 -45 1070
rect 35 1045 55 1130
rect -25 1035 55 1045
rect -25 1015 -15 1035
rect 5 1025 55 1035
rect 5 1015 15 1025
rect -25 1005 15 1015
rect -65 965 15 985
rect -5 770 15 965
rect 75 895 95 1170
rect 115 945 155 955
rect 115 925 125 945
rect 145 935 155 945
rect 145 925 175 935
rect 115 915 175 925
rect 75 875 115 895
rect 95 865 135 875
rect 95 845 105 865
rect 125 845 135 865
rect 95 835 135 845
rect 155 810 175 915
rect 95 790 175 810
rect 95 770 115 790
rect -110 760 -70 770
rect -110 690 -100 760
rect -80 690 -70 760
rect -110 680 -70 690
rect -5 760 35 770
rect -5 690 5 760
rect 25 690 35 760
rect -5 680 35 690
rect 75 760 115 770
rect 75 690 85 760
rect 105 690 115 760
rect 75 680 115 690
rect 140 760 180 770
rect 140 690 150 760
rect 170 690 180 760
rect 140 680 180 690
rect -35 630 5 640
rect -35 560 -25 630
rect -5 560 5 630
rect -35 550 5 560
rect 100 630 140 640
rect 100 560 110 630
rect 130 560 140 630
rect 100 550 140 560
rect -115 520 185 530
rect -115 510 -80 520
rect -90 500 -80 510
rect -60 510 40 520
rect -60 500 -50 510
rect -90 490 -50 500
rect 30 500 40 510
rect 60 510 185 520
rect 60 500 70 510
rect 30 490 70 500
<< viali >>
rect -45 2060 -25 2130
rect 95 2060 115 2130
rect 30 1905 50 1975
rect 30 1375 50 1445
rect -100 1180 -80 1250
rect 150 1180 170 1250
rect -100 690 -80 760
rect 150 690 170 760
rect -25 560 -5 630
rect 110 560 130 630
<< metal1 >>
rect -135 2130 205 2165
rect -135 2060 -45 2130
rect -25 2060 95 2130
rect 115 2060 205 2130
rect -135 2025 205 2060
rect 20 1975 60 2025
rect 20 1905 30 1975
rect 50 1905 60 1975
rect 20 1445 60 1905
rect 20 1375 30 1445
rect 50 1375 60 1445
rect 20 1365 60 1375
rect -115 1250 -70 1265
rect -115 1180 -100 1250
rect -80 1180 -70 1250
rect -115 760 -70 1180
rect -115 690 -100 760
rect -80 690 -70 760
rect -115 645 -70 690
rect 140 1250 185 1265
rect 140 1180 150 1250
rect 170 1180 185 1250
rect 140 760 185 1180
rect 140 690 150 760
rect 170 690 185 760
rect 140 645 185 690
rect -115 630 185 645
rect -115 560 -25 630
rect -5 560 110 630
rect 130 560 185 630
rect -115 545 185 560
<< labels >>
rlabel locali -115 520 -115 520 7 CLK
port 1 w
rlabel metal1 -135 2095 -135 2095 7 VDD
port 2 w
rlabel metal1 -115 595 -115 595 7 GND
port 3 w
rlabel pdiff -115 1940 -115 1940 7 D
port 4 w
rlabel pdiff -115 1410 -115 1410 7 Dn
port 5 w
rlabel pdiff 185 1940 185 1940 3 Q
port 6 e
rlabel locali 180 1410 180 1410 3 Qn
port 7 e
<< end >>
